** Profile: "SCHEMATIC1-last run of dc sweep "  [ D:\A\e, sources\Electrical Circuit\Project\Final project _1\Final Project-SCHEMATIC1-last run of dc sweep .sim ] 

** Creating circuit file "Final Project-SCHEMATIC1-last run of dc sweep .sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\..\..\..\..\orcad\capture\library\pspice\Final Project-SCHEMATIC1.net" 


.END
