** Profile: "SCHEMATIC1-last run"  [ D:\A\e, sources\Electrical Circuit\Homeworks\hw9\9431022-yasaman mirmohammad-hw9\4\9-4-SCHEMATIC1-last run.sim ] 

** Creating circuit file "9-4-SCHEMATIC1-last run.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\9-4-SCHEMATIC1.net" 


.END
