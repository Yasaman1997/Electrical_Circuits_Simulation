** Profile: "SCHEMATIC1-5th run"  [ D:\A\e, sources\Electrical Circuit\Homeworks\hw8\1\8-1-SCHEMATIC1-5th run.sim ] 

** Creating circuit file "8-1-SCHEMATIC1-5th run.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\8-1-SCHEMATIC1.net" 


.END
