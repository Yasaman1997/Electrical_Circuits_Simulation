** Profile: "SCHEMATIC1-4-b"  [ D:\A\e, sources\Electrical Circuit\Homeworks\hw8\4\8-4-schematic1-4-b.sim ] 

** Creating circuit file "8-4-schematic1-4-b.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC DEC PARAM a 100 100k 20 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\8-4-SCHEMATIC1.net" 


.END
