** Profile: "SCHEMATIC1-last run"  [ D:\A\e, sources\Electrical Circuit\Project\Final project _1\Final Project-SCHEMATIC1-last run.sim ] 

** Creating circuit file "Final Project-SCHEMATIC1-last run.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 1 1 meg 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\..\..\..\..\orcad\capture\library\pspice\Final Project-SCHEMATIC1.net" 


.END
