** Profile: "SCHEMATIC1-last dc sweep run"  [ D:\A\e, sources\Electrical Circuit\Project\Final project _1\final project-schematic1-last dc sweep run.sim ] 

** Creating circuit file "final project-schematic1-last dc sweep run.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM a 0.5 4 0.001 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\..\..\..\..\orcad\capture\library\pspice\Final Project-SCHEMATIC1.net" 


.END
